class frame_info_struct extends uvm_component;
endclass
